module practica_minios (clock, reset, LEDS);

input clock;
input reset;
output [7:0] LEDS;


endmodule