
module DE0_NANO_SOPC (
	clk_clk,
	pio_led_external_connection_export);	

	input		clk_clk;
	output	[7:0]	pio_led_external_connection_export;
endmodule
